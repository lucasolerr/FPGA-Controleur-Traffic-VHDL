Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;


entity constante7 is
PORT (
		sept: out std_logic_vector (2 downto 0)
		

		
);
end constante7;

architecture DESCRIPTION of constante7 is

begin

	
	sept <= "111"; --7

end DESCRIPTION;